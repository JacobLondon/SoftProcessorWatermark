`timescale 1ns / 1ps

module RegisterFile(
    write,
    address1,
    address2,
    address3,
    valRead1,
    valRead2,
    valWrite3,
    clk
);

input readwrite;            // read == 0, write == 1
input [4:0] address1;       // read: address of register 1
input [4:0] address2;       // read: address of register 2

output [31:0] valRead1;     // read: value of register 1
output [31:0] valRead2;     // read: value of register 2

input [4:0] address3;       // write: address of register 3
input [31:0] valWrite3;     // write: value of register 3

input clk;

// initialize register memory
reg [31:0] rmemory [31:0];

// table generated by format.py
initial begin
    
    rmemory[0] = 32'b00000000000000000000000000000000;
    rmemory[1] = 32'b00000000000000000000000000000000;
    rmemory[2] = 32'b00000000000000000000000000000000;
    rmemory[3] = 32'b00000000000000000000000000000000;
    rmemory[4] = 32'b00000000000000000000000000000000;
    rmemory[5] = 32'b00000000000000000000000000000000;
    rmemory[6] = 32'b00000000000000000000000000000000;
    rmemory[7] = 32'b00000000000000000000000000000000;
    rmemory[8] = 32'b00000000000000000000000000000000;
    rmemory[9] = 32'b00000000000000000000000000000000;
    rmemory[10] = 32'b00000000000000000000000000000000;
    rmemory[11] = 32'b00000000000000000000000000000000;
    rmemory[12] = 32'b00000000000000000000000000000000;
    rmemory[13] = 32'b00000000000000000000000000000000;
    rmemory[14] = 32'b00000000000000000000000000000000;
    rmemory[15] = 32'b00000000000000000000000000000000;
    rmemory[16] = 32'b00000000000000000000000000000000;
    rmemory[17] = 32'b00000000000000000000000000000000;
    rmemory[18] = 32'b00000000000000000000000000000000;
    rmemory[19] = 32'b00000000000000000000000000000000;
    rmemory[20] = 32'b00000000000000000000000000000000;
    rmemory[21] = 32'b00000000000000000000000000000000;
    rmemory[22] = 32'b00000000000000000000000000000000;
    rmemory[23] = 32'b00000000000000000000000000000000;
    rmemory[24] = 32'b00000000000000000000000000000000;
    rmemory[25] = 32'b00000000000000000000000000000000;
    rmemory[26] = 32'b00000000000000000000000000000000;
    rmemory[27] = 32'b00000000000000000000000000000000;
    rmemory[28] = 32'b00000000000000000000000000000000;
    rmemory[29] = 32'b00000000000000000000000000000000;
    rmemory[30] = 32'b00000000000000000000000000000000;
    rmemory[31] = 32'b00000000000000000000000000000000;

end

// read
assign valRead1 = rmemory[address1];
assign valRead2 = rmemory[address2];

// write
always @(negedge clk) begin
    // if writing
    if(readwrite==1'b1) begin
        rmemory[address3] = valWrite3;
    end
end

endmodule