`timescale 1ns / 1ps

module InstructionMemory(inst, pc, clk);
input clk;
input  [31:0] pc;
output [31:0] inst;
reg    [31:0] inst;

// initialize inst memory
reg [31:0] memdata [127:0];


// generate insts here
// http://www.kurtm.net/mipsasm
initial begin

// test program
/*
    memdata[0] = 32'b00000001110011100111000000100010;
    memdata[1] = 32'b00000000000011001000001000000010;
    memdata[2] = 32'b00000000000011011000101000000010;
    memdata[3] = 32'b00000010000100011010100000100000;
    memdata[4] = 32'b00000000000101011010100001000010;
    memdata[5] = 32'b00000000000101011010101000000000;
    memdata[6] = 32'b00000001110101010111000000100101;
    memdata[7] = 32'b00000001100100111000000000100100;
    memdata[8] = 32'b00000000000100001000000100000010;
    memdata[9] = 32'b00000001101100111000100000100100;
    memdata[10] = 32'b00000000000100011000100100000010;
    memdata[11] = 32'b00000010000100011010100000100000;
    memdata[12] = 32'b00000000000101011010100001000010;
    memdata[13] = 32'b00000000000101011010100100000000;
    memdata[14] = 32'b00000001110101010111000000100101;
    memdata[15] = 32'b00000001100101001000000000100100;
    memdata[16] = 32'b00000001101101001000100000100100;
    memdata[17] = 32'b00000010000100011010100000100000;
    memdata[18] = 32'b00000000000101011010100001000010;
    memdata[19] = 32'b00000001110101010111000000100101;
    memdata[20] = 32'b00000000000000000000000000000000;

*/
    // nothing
    //memdata[0] = 32'b00000000000000000000000000000000;

    // program
    memdata[0] = 32'b00000001110011100111000000100010;
    memdata[1] = 32'b00000000000011001000001000000010;
    memdata[2] = 32'b00000000000011011000101000000010;
    memdata[3] = 32'b00000010000100011010100000100000;
    memdata[4] = 32'b00000000000101011010100001000010;
    memdata[5] = 32'b00000000000101011010101000000000;
    memdata[6] = 32'b00000001110101010111000000100101;
    memdata[7] = 32'b00000001100100111000000000100100;
    memdata[8] = 32'b00000000000100001000000100000010;
    memdata[9] = 32'b00000001101100111000100000100100;
    memdata[10] = 32'b00000000000100011000100100000010;
    memdata[11] = 32'b00000010000100011010100000100000;
    memdata[12] = 32'b00000000000101011010100001000010;
    memdata[13] = 32'b00000000000101011010100100000000;
    memdata[14] = 32'b00000001110101010111000000100101;
    memdata[15] = 32'b00000001100101001000000000100100;
    memdata[16] = 32'b00000001101101001000100000100100;
    memdata[17] = 32'b00000010000100011010100000100000;
    memdata[18] = 32'b00000000000101011010100001000010;
    memdata[19] = 32'b00000001110101010111000000100101;
    memdata[20] = 32'b00000001011010010101100000100000; // add counter
    memdata[21] = 32'b00010001011010100000000000000001; // beq 1
    memdata[22] = 32'b00010101000010011111111111101001; // bne -23
    memdata[23] = 32'b00000001011010110101100000100010; // sub
    memdata[24] = 32'b00010101000010011111111111100111; // bne -25
    memdata[25] = 32'b00000000000000000000000000000000;

end

// set the next inst
always @(posedge clk) begin
    inst = memdata[pc];
end

endmodule
